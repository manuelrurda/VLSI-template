LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY practica1 IS
	PORT ()
	

END practica1;

ARCHITECTURE BEHAVIORAL OF practica1 IS
	
	BEGIN
	
	
	
END ARCHITECTURE;
