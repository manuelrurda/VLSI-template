"00010001" --A
"00000001"--B
"01100011"--C
"10000101"--D
"01100001"--E
"01110001"--F
"01000001"--G
"10010001"--H
"10011111"--I
"10000111"--J
"10010001"--K
"10011101"--L
"11010101"--M
"11010101"--N
"00000011"--O
"00110001"--P
"00110001"--Q
"00010001"--R
"01001001"--S
"11100001"--T
"10000011"--U
"10000011"--V
"10010001"--W
"10010001"--X
"10011001"--Y
"00100101"--Z
"00010001"--a
"11000001"--b
"11100101"--c
"10000101"--d
"01100001"--e
"01110001"--f
"00001001"--g
"11010001"--h
"11011111"--i
"10001111"--j
"10010001"--k
"10011111"--l
"11010101"--m
"11010101"--n
"00000011"--o
"00110001"--p
"00110001"--q
"11110101"--r
"01001001"--s
"11100001"--t
"11000111"--u
"11000111"--v
"00000001"--w
"10010001"--x
"10011001"--y
"00100101"--z
"00000011"--0
"10011111"--1
"00100101"--2
"00001101"--3
"10011001"--4
"01001001"--5
"01000001"--6
"00011111"--7
"00000001"--8
"00110001"--9
--ABCDEFG.
  
